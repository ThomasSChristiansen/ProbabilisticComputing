`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT(group_EN, Pbit_EN);

input logic [0:2] group_EN;
output logic [0:222] Pbit_EN;

always_comb
begin 
case (group_EN)
  3'b000 : Pbit_EN = 223'b0010000100100100010001001000010000000101000010101001001001001001001001000100010010000101000100001010000010100000000100000100000010000010100000000001010001001010000010000000101000100101000000000100010111111010000000000101111;
  3'b001 : Pbit_EN = 223'b0000001001001000001000100110100110001000101001000010000010000000000000001001000100100000010001000001001000010010010010010000010100000101001000100010100000100100110100010001010000010000001001100001000000000001011011001010000;
  3'b010 : Pbit_EN = 223'b0100010000010010100100010001000001010000010100000000010000100010010010010010001000010010001000100100010001000100100000100010001000010000010101011000000100000000000001001100000010001000010100010000001000000000100100110000000;
  3'b011 : Pbit_EN = 223'b1001100010000001000010000000001000100010000000010100100100010100100100100000100001001000100010010000100100001001001001001001100001101000000010000100001010010001001000100010000101000010100010001010100000000100000000000000000;
endcase
end
endmodule
