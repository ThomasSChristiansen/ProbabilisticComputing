`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT(group_EN, Pbit_EN);

input logic [0:2] group_EN;
output logic [0:458] Pbit_EN;

always_comb
begin 
case (group_EN)
  3'b000 : Pbit_EN = 459'b010001000100001001001001000010010010000001001000000001010001010001010000100010000000101000000010001000001010001000100001001000100100000001000100000010000100010001000100100100010010010000010001000100000100100100100100000100100100101000100010000001001000010100001000000110001010000001011000010001000101000000001000000000100100010011000001100000100001000000000110010000000000000000000010100010100100001000000010100010100010000000011111111000000000011111110110111;
  3'b001 : Pbit_EN = 459'b000010010000010010010010000101000100100010010010110000000100000100000100000100101010000010001000010110100000000100001000100100010000010100100000100000100011100000100000001001000100100010001010000011001010010001000000100001010000010100010001000010000101100001000000100000100001110010000010000000010000010010100111100000010010000000001000001000001000010001001001000100110000001001110000000001001011010001110000000000010000101000100000000010101101100000001001000;
  3'b010 : Pbit_EN = 459'b000100000011100000000000101000101000011100000001001110001000100000100001010000010100010001100100000000010001010001000100000010000001001010001001011000000000000100001001000000100001001000100100010000110000001000001010001000001010000010000100111000100000000010010011010001000100001000000101100100100010000100010000010101000000101000010010010010000010001100100000001010001000000110000101001000000000000100000101001001001001010001000000000101010010000000000000000;
  3'b011 : Pbit_EN = 459'b101000101000000100100100010000000001000000100100000000100010001010001010001001000001000100010001000001000100100010010010010001001010100000010010000101001000001010010010010010001000000101000000101000000001000010010001010010000001000001001000000100010010001000100100001000010000000100100000001010001000101001000000001010001001000100100100000101010100100010010000100001000111110000001000010100010000100010001000010100000100000110000000000000000000000000000000000;
  3'b100 : Pbit_EN = 459'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule
