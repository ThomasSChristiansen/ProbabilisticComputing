`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT(group_EN, Pbit_EN);

input logic [0:2] group_EN;
output logic [0:993] Pbit_EN;

always_comb
begin 
case (group_EN)
  3'b000 : Pbit_EN = 994'b0101000100000000100100000001010001010001000100010000010000000101000000010100010100010010100010000010000010001000100000010010010000000010001001000001001001000001010010010000001000001000001010001000100100100100000010010001000010001000010001010000100001000001000001010001000100100000100100010010001001000100001010000100100100001000001000010000010100010001001000001000001001001000100110001001000010001100000100100010000100000000100100001100100010000100100000000000000000101000100110000001001000010100001001001000011001001001000100001001000000010010000101000100000001000000100000100010011010000010000001000100010100010010010010001001000001010000001100100000001001000101000010100010000000100010010000010000100000101010000001000100010100000101000001001001000001010000001000100000010001000101000100010100001001000001010010001000010000100000100010010001001000001001000001000100100010001001000001000010010101001001000100001001010001001001000110000000000000111111101111111100000000000000000000111110110100;
  3'b001 : Pbit_EN = 994'b0010000001001001001001100010100000000000100010001011000110001010010000101001000000000000000100000101110100100000010010000100000010100001000000001000100010101000100100000101000100010100010100000100000001000001001000000010010100010101000100000100001000100010100010100000100000001001000001001001000000010001000101010001000001000010010000101000101000001000000010010001000100010001001000100010010000010010010001001001000001001010001010010001000001000000001001011000101000010010000000010100010010001001000010010101000010010000000010010010101100100100000000000001001000001100000100000001000101100100010100001000001001100000001100100010010100000110010001001100100010000000000000000000100100000100001001001100011001000100110000100010000001100000011100000100101000000110010100010100101000100010000000000000100000001000100100010001000110001001001000001010000010100000010010001001001000010000100010101000000000100000001010010010001000000000010000100100010000000000000000000010111001110101100111000001001011;
  3'b010 : Pbit_EN = 994'b0000101010100110000000011000000100100100010001000000100001100000001010000010001001001001010001010000001000000101001001000000100101001000010100010100000100000110001000100010100010000011000000100001001000001000100101001000000001000010100000100010010100010000011000000100001001000100001010000000010010101000100000101000001000100101000100000110000001000010010001000010010000100100000000010000100101000001101000000100010010100100000001100000001000011001000100100010010010000001001000101010000001000000100000000010100000000010110001100000000011000001010010010010010010100001010001011000000000010001001010000001000010000101000001010000001000100001100000000011000000010010101001001000001010001001000010000001000010000001001010000001001000010010000010010000010000100001000010001010000100010000001001001001000100100100000001000110100001000010000100100000010001010010001100100000000100000100001100010001001000000100100001100000000100100100000000010011001000000000010000000001000110001010011000000000000000;
  3'b011 : Pbit_EN = 994'b1000010000010000010010000100001010001010001000100100001000010000100101000000100010100100001000101000000001010010000100001001001000010100100010100010010000010000000001001000010001000000100001010010010010010010010000100100101000100000001010001001000010001000000100001010010010010010010000100100100100000010010000000010010010010000100010000001000010100100100100100100100010000010010001000100001000100000000010010000101000010000010000000010010100100010010010000101000101000100010001000000100100100010010100100000000100100100001000000100010000001000101000101000100100010010001010000100100000001000100000110010100000001000100000000100100010001000000010010000010100101000010100010101010001010000100100100010000100010000000100011000100010001000100000100010000110001000100001000001000010001000110010100010010010010010001000100000001000010100010001000100100100000100100000010010010001100010010000000100100010010010010000000100100010010010101001001000100111000000000000000000000000000000000000000000000000;
  3'b100 : Pbit_EN = 994'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule
