`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT(group_EN, Pbit_EN);

input logic [0:2] group_EN;
output logic [0:45] Pbit_EN;

always_comb
begin 
case (group_EN)
  3'b000 : Pbit_EN = 46'b0110000000100100101000100100000100101000000111;
  3'b001 : Pbit_EN = 46'b0001010001000000010001010000100010000011000000;
  3'b010 : Pbit_EN = 46'b1000001010001010000100000010010000010100011000;
  3'b011 : Pbit_EN = 46'b0000100100010001000010001001001001000000100000;
endcase
end
endmodule
