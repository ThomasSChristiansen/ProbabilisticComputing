// pbit_params.svh
// Global parameter definitions for all p-bit modules

`ifndef GLOBAL_PARAMS_SVH
`define GLOBAL_PARAMS_SVH

// Define the number of P-bits globally
parameter num_Pbits = 46;
parameter num_Out = 
parameter HIST_DATA_SIZE = 63;`endif
