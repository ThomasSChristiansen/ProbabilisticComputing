// pbit_params.svh
// Global parameter definitions for all p-bit modules

`ifndef GLOBAL_PARAMS_SVH
`define GLOBAL_PARAMS_SVH

// Define the number of P-bits globally
parameter num_Pbits = 994;

`endif
