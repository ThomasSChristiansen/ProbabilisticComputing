`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT(group_EN, Pbit_EN);

input logic [0:2] group_EN;
output logic [0:90] Pbit_EN;

always_comb
begin 
case (group_EN)
  3'b000 : Pbit_EN = 91'b0001000110010000000001000100100010101100000010000010011001000000000100010001101000000111110;
  3'b001 : Pbit_EN = 91'b0110010000000100111000001000001001010000010000010000000010001001010001000000010000001000001;
  3'b010 : Pbit_EN = 91'b0000100001001010000100010001000100000001000100101000100000100100100010001000000111100000000;
  3'b011 : Pbit_EN = 91'b1000001000100001000010100010010000000010101001000101000100010010001000100110000000010000000;
endcase
end
endmodule
