`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT(group_EN, Pbit_EN);

input logic [0:2] group_EN;
output logic [0:2022] Pbit_EN;

always_comb
begin 
case (group_EN)
  3'b000 : Pbit_EN = 2023'b0000101000100010010000000000010000100000010001000000100110001010000010100000000100100001001000000010010000010000101000101000010100010010001001011000100000000100010001000100100000001001000010100001010000000010010100010100000001001001100100100100010010010001001001000100110100011000101000001001000000010010001001000010100010000100100000101000000010010001001000010000001000001000000000110110001000100100001001000000010010000101000011010000000100010000101000001000100010100001000000100000000010000010000100000011001000000010010001011000010100000000100100000100100000010010010011001000001000000001001010001010000010010000000100100010010010010011000010010000101000000001000001000100100011100101001000100000000100010000001000100010100000100100001000100010000010001000000100110000010010010000010010001000010010000101000010001000100000010000100000000110001010010010011000010010000000100100001010000100010000000010001000100011100100100010000100100000010001001000100000000000001000111000010101000010010001001000010100000000000011100010010000001000100010010110000000000010000001010100100000000100100000011101000000010000000100010100100000001001001000100000010001000100001000010010010001000010001000000001000001000100100001000100000101000000010100010100010000000001000100010100010010000000100100001010000000101000000010100010100010100010100000100100100011000000100001000000100010001010000001001000000010100010100010100010100010001001000100000000101000010001000000101000010100000001010000000101000101000101000100010000010010001001000000010100010100010001000000010100001010000000101000000010100010100001010001010000100100001001001000000001000001001010001001000010100000000100100000101000010001010000000010100010010001010010101000101000100100000000010000001001000000010010001010000010100000000100100000101000000001010000000001010001101000101000010100010000100000100101000001010000000010001000000100010001010001010100000000100100001101000000010010000000100100010100101010001011111111111111111000000000000000000101101110011110111111101111111;
  3'b001 : Pbit_EN = 2023'b0000000000010100100100001101000100011111000000011110000000000000101000001111100000001000100011110001000111100010000000000000000000000000000000100010011110010001001110110000001001100000010000001000000011111000000010000001111100000010000000000000000000000000000000000000001001000010010111100000011111000000000000010000001101110000000100000011110001000000100010000011000001000000100100001000100010010011100000001111000000000000010000000111110010000100000001110000001000001000010100000100010001101000001001111000000011110000000000000010000001101100000001100000000100000000000100000001000010100100010000010001101000000111010000000000000100000000110001000100010000100010100010100000001000001000010001001001110000000111100000000000000100000011100000010000110100010101010000000000100000101011000000110110000000010000010000000001010011000101001010110000100000100000100111000000101100010000000000100000000010010001000010000100001000001101110000010111100000100000010010001001000100000010000010111000000010000001000010010001000100001000100111000100000000001000100100100001101000001011001001000000000101000000000100100100100010001000010001010000010101001111000100000011100000000000000100001000010001001000001010110000001000100011100000011110000000000000001001001000001011000001001000111110000001000000111100000011110000000000000000000000001000000000011000011010000100111110000001000000111100000011110000000000000000000000000001000100100000111100000010001000111100000010000001111000000111100000000000000000000010000010000000010010111110000000000001000100111110000001000000111100000011110000000000000000000000000000010010000010000111010000101110000000000110010000001111110000000100000011101000000111010000000000000000000000000000000000001001001110001111000000011110000000000001010000001111110000001100000011111000000111100000000000000000000000000000001000000100001000101000100011111000000011110000000000000100000001111100000001000000011110000000111010010000000000000000000000000000000000000010010010010010110010010001100001000000010000000;
  3'b010 : Pbit_EN = 2023'b0101000101000000001001110010100000000000100110000001001000100100010001000000001001000100010000000000100000000100010010010001001001001100100100000000000001101000000000001001000100010010000101000100100000000100100001001000000010100100001001010010101000101000010100011001000010100000000000010010000000100100100110001001000000001001000001000100000100001010000100101000010100010011010001000001010000000000010010010000100100010010000100001000000000100001000110000010010001000010100001010010001000010001100010000100010000001100100100100000100010000011010010001010001010001000100000010100010100010010100001000100000100100000101001001000100000101000000100001001000010010000001000010010010100000010100010000010001010100000000001001001001001010000010010000100001001000000100010000111000100000000100100000001101001001000100101100010000100000010000100001001010101000100000000100100000001000010110001001010001001000100100001001000010001000000000001000000000100010010000100010100010010000100100000000101001100010010001000100100010000010001000000010000010100100000001001001100010010000000000010010010001000100010000001000001001000100010001100000010000000000000100000101000010010000100101010010001000010100100010100001001000100001000001010000000101001001001000010010100010000000000100001000001001000100100000001010000000101001001001001001001000010010010000000100101001000000001001000100100000010010000000101001001001001001001001000100010001001000001010000100010000001010001001000000010100000001010010010010010010000100100101000100000000000101001001000100000000000101000100100000001010000000101001001001100100100100010000001010000100000101010000000010100100000101001000000001001001010010000000010100000000001001001100100100100010010010001000000010001000000110010000001000100100100001001000000001001000010010000000010100000011110001010000101000100100010100011001010000010010100000000000100110000001001000100100010001000000011001000100010000000100100000001000010100010010001010000000000000000000101101101101101001000000000000000000000000000000;
  3'b011 : Pbit_EN = 2023'b1010010010001001000010000000001011000000001000100000010001010001000100010000010010010010000100001100001000001001000101000110100010100001010010000101000000000010100000000010010010000100101000010010001100000001001000100010000000010000010010001001000101000110100010100010000000000101000000000100100000001001010000100100010000000010011010010000001000100100010001000100100010100100001010000000000101001000000100100000001001101000101000100000001001001010010000000101000100010100001010001001100100000100010000000000100100000001001010000101001000010000001000010001010001100101001000100010100001001000000100100000010001001000000010010101001001000100001000100010000101001100010100001001000000010000000100000100000001001000010110010100010010001000000101001001000000100010001001001000001001000100001001000000000100100010001000010100001000101000010001000000000000001001000000001001010010001001000100010001100100101000010100010000000010010000001010001000001010000101001001100010100001000001001000000000100000100100100001001010101000000100001000100011001001000001010010010000000100100000010100101001010010000000111010001010010001000001000010100100100010010000001010010000000100101001000000100100100100010010100000000010010010010000010000100001000010100010100100100010100000101010000100000000010010010001000010000100001000010100010100010100010101001001000100000000010010000000010100010001000000100100001000010100010100010100010100010000010010000010000101000100000010000100100010000100001000010000101000101000101001001001000101000100000001000010100010001010000001000010010001000010000100001000010100010010001010001101001000100100010000000100010000100001010000000100010000000010010001000100000100001000101100010100001010001001000101000110010010100000100000000100100000101001010000100100010000000010010001000100000100001000000000100100010010010011001001000100010001010000000010001100000001000100000010101010001000100010000000010010010000100001001001000100001001001001000100100100000000000000000000000000000000000000000000000000000000000000000;
  3'b100 : Pbit_EN = 2023'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
endcase
end
endmodule
