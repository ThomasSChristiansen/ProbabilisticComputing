`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////


module grouped_update_order_LUT #(
    parameter num_Pbits = 4
)(
    input logic [0:3] group_EN,
    output logic [0:num_Pbits-1] Pbit_EN
);

always_comb
begin 
case (group_EN)
3'b000 : Pbit_EN = 53'b11110000000000000000000000001010000000010100000001011;
3'b001 : Pbit_EN = 53'b00001011011000000100000000110100000000001000000000100;
3'b010 : Pbit_EN = 53'b00000100000100000000101000000001010000100000101100000;
3'b011 : Pbit_EN = 53'b00000000100000010000000111000000000111000010010010000;
3'b100 : Pbit_EN = 53'b00000000000011101011010000000000101000000001000000000;
endcase
end
endmodule